
/////////////////////// Testbench for B2T///////////////////

module tb_bin_to_thermo;

// Testbench signals
reg  [3:0] binary;
wire [15:0] thermo;
// Instantiate the bin_to_thermo module
B2T uut (
	.binary(binary),
	.thermo(thermo)
);
initial begin
	// Display signal values on each change
  $monitor("Time = %0d, binary = %b, decimal = %d, thermo = %b", $time, binary,binary, thermo);
	// Test all binary input values
	binary = 4'b0000; #10;
	binary = 4'b0001; #10;
	binary = 4'b0010; #10;
	binary = 4'b0011; #10;
	binary = 4'b0100; #10;
	binary = 4'b0101; #10;
	binary = 4'b0110; #10;
	binary = 4'b0111; #10;
	binary = 4'b1000; #10;
	binary = 4'b1001; #10;
	binary = 4'b1010; #10;
	binary = 4'b1011; #10;
	binary = 4'b1100; #10;
	binary = 4'b1101; #10;
	binary = 4'b1110; #10;
	binary = 4'b1111; #10;
	// Finish the simulation
	$finish;
end
endmodule



